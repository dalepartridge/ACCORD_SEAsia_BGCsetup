netcdf nemoersem_ini_trc {
dimensions:
	y = 375 ;
	x = 297 ;
	z = 51 ;
	t = UNLIMITED ; // (1 currently)
variables:
	double kt ;
		kt:long_name = "number of time steps" ;
		kt:units = "1" ;
	double time_counter(t) ;
		time_counter:long_name = "number of time steps" ;
		time_counter:units = "1" ;
	double rdttrc1 ;
		rdttrc1:long_name = "time step" ;
		rdttrc1:units = "s" ;
	float nav_lat(y, x) ;
		nav_lat:long_name = "latitude" ;
		nav_lat:units = "degrees_north" ;
	float nav_lon(y, x) ;
		nav_lon:long_name = "longitude" ;
		nav_lon:units = "degrees_east" ;
	float nav_lev(z) ;
		nav_lev:long_name = "vertical levels" ;
		nav_lev:units = "1" ;
	double adatrj ;
		adatrj:long_name = "days since the beginning of the run" ;
		adatrj:units = "d" ;
	double TRNP1_c(t, z, y, x) ;
		TRNP1_c:long_name = "diatom carbon" ;
		TRNP1_c:units = "mg/m3" ;
	double TRNP1_n(t, z, y, x) ;
		TRNP1_n:long_name = "diatom nitrogen" ;
		TRNP1_n:units = "mmol/m3" ;
	double TRNP1_p(t, z, y, x) ;
		TRNP1_p:long_name = "diatom phosphate" ;
		TRNP1_p:units = "mmol/m3" ;
	double TRNP1_s(t, z, y, x) ;
		TRNP1_s:long_name = "diatom silicate" ;
		TRNP1_s:units = "mmol/m3" ;
	double TRNP1_Chl(t, z, y, x) ;
		TRNP1_Chl:long_name = "diatom chlorophyll-a" ;
		TRNP1_Chl:units = "mg/m3" ;
	double TRNP2_c(t, z, y, x) ;
		TRNP2_c:long_name = "nanophytoplankton carbon" ;
		TRNP2_c:units = "mg/m3" ;
	double TRNP2_n(t, z, y, x) ;
		TRNP2_n:long_name = "nanophytoplankton nitrogen" ;
		TRNP2_n:units = "mmol/m3" ;
	double TRNP2_p(t, z, y, x) ;
		TRNP2_p:long_name = "nanophytoplankton phosphate" ;
		TRNP2_p:units = "mmol/m3" ;
	double TRNP2_Chl(t, z, y, x) ;
		TRNP2_Chl:long_name = "nanophytoplankton chlorophyll-a" ;
		TRNP2_Chl:units = "mg/m3" ;
	double TRNP3_c(t, z, y, x) ;
		TRNP3_c:long_name = "picophytoplankton carbon" ;
		TRNP3_c:units = "mg/m3" ;
	double TRNP3_n(t, z, y, x) ;
		TRNP3_n:long_name = "picophytoplankton nitrogen" ;
		TRNP3_n:units = "mmol/m3" ;
	double TRNP3_p(t, z, y, x) ;
		TRNP3_p:long_name = "picophytoplankton phosphate" ;
		TRNP3_p:units = "mmol/m3" ;
	double TRNP3_Chl(t, z, y, x) ;
		TRNP3_Chl:long_name = "picophytoplankton chlorophyll-a" ;
		TRNP3_Chl:units = "mg/m3" ;
	double TRNP4_c(t, z, y, x) ;
		TRNP4_c:long_name = "microphytoplankton carbon" ;
		TRNP4_c:units = "mg/m3" ;
	double TRNP4_n(t, z, y, x) ;
		TRNP4_n:long_name = "microphytoplankton nitrogen" ;
		TRNP4_n:units = "mmol/m3" ;
	double TRNP4_p(t, z, y, x) ;
		TRNP4_p:long_name = "microphytoplankton phosphate" ;
		TRNP4_p:units = "mmol/m3" ;
	double TRNP4_Chl(t, z, y, x) ;
		TRNP4_Chl:long_name = "microphytoplankton chlorophyll-a" ;
		TRNP4_Chl:units = "mg/m3" ;
	double TRNZ4_c(t, z, y, x) ;
		TRNZ4_c:long_name = "mesozooplankton carbon" ;
		TRNZ4_c:units = "mg/m3" ;
	double TRNZ5_c(t, z, y, x) ;
		TRNZ5_c:long_name = "microzooplankton carbon" ;
		TRNZ5_c:units = "mg/m3" ;
	double TRNZ5_n(t, z, y, x) ;
		TRNZ5_n:long_name = "microzooplankton nitrogen" ;
		TRNZ5_n:units = "mmol/m3" ;
	double TRNZ5_p(t, z, y, x) ;
		TRNZ5_p:long_name = "microzooplankton phosphorus" ;
		TRNZ5_p:units = "mmol/m3" ;
	double TRNZ6_c(t, z, y, x) ;
		TRNZ6_c:long_name = "heteroflagellates carbon" ;
		TRNZ6_c:units = "mg/m3" ;
	double TRNZ6_n(t, z, y, x) ;
		TRNZ6_n:long_name = "heteroflagellates nitrogen" ;
		TRNZ6_n:units = "mmol/m3" ;
	double TRNZ6_p(t, z, y, x) ;
		TRNZ6_p:long_name = "heteroflagellates phosphorus" ;
		TRNZ6_p:units = "mmol/m3" ;
	double TRNB1_c(t, z, y, x) ;
		TRNB1_c:long_name = "particualte organic carbon" ;
		TRNB1_c:units = "mg/m3" ;
	double TRNB1_n(t, z, y, x) ;
		TRNB1_n:long_name = "particualte organic nitrogen" ;
		TRNB1_n:units = "mmol/m3" ;
	double TRNB1_p(t, z, y, x) ;
		TRNB1_p:long_name = "particualte organic phosphorus" ;
		TRNB1_p:units = "mmol/m3" ;
	double TRNR1_c(t, z, y, x) ;
		TRNR1_c:long_name = "dissolved organic carbon" ;
		TRNR1_c:units = "mg/m3" ;
	double TRNR1_n(t, z, y, x) ;
		TRNR1_n:long_name = "dissolved organic nitrogen" ;
		TRNR1_n:units = "mmol/m3" ;
	double TRNR1_p(t, z, y, x) ;
		TRNR1_p:long_name = "dissolved organic phosphorus" ;
		TRNR1_p:units = "mmol/m3" ;
	double TRNR2_c(t, z, y, x) ;
		TRNR2_c:long_name = "semi-labile organic carbon" ;
		TRNR2_c:units = "mg/m3" ;
	double TRNR3_c(t, z, y, x) ;
		TRNR3_c:long_name = "semi-refractory organic carbon" ;
		TRNR3_c:units = "mg/m3" ;
	double TRNR4_c(t, z, y, x) ;
		TRNR4_c:long_name = "small particulate organic carbon" ;
		TRNR4_c:units = "mg/m3" ;
	double TRNR4_n(t, z, y, x) ;
		TRNR4_n:long_name = "small particulate organic nitrogen" ;
		TRNR4_n:units = "mmol/m3" ;
	double TRNR4_p(t, z, y, x) ;
		TRNR4_p:long_name = "small particulate organic phosphorus" ;
		TRNR4_p:units = "mmol/m3" ;
	double TRNR6_c(t, z, y, x) ;
		TRNR6_c:long_name = "medium size particulate organic carbon" ;
		TRNR6_c:units = "mg/m3" ;
	double TRNR6_n(t, z, y, x) ;
		TRNR6_n:long_name = "medium size particulate organic nitrogen" ;
		TRNR6_n:units = "mmol/m3" ;
	double TRNR6_p(t, z, y, x) ;
		TRNR6_p:long_name = "medium size particulate organic phosphorus" ;
		TRNR6_p:units = "mmol/m3" ;
	double TRNR6_s(t, z, y, x) ;
		TRNR6_s:long_name = "medium size particulate organic silicate" ;
		TRNR6_s:units = "mmol/m3" ;
	double TRNR8_c(t, z, y, x) ;
		TRNR8_c:long_name = "large particulate organic carbon" ;
		TRNR8_c:units = "mg/m3" ;
	double TRNR8_n(t, z, y, x) ;
		TRNR8_n:long_name = "large particulate organic nitrogen" ;
		TRNR8_n:units = "mmol/m3" ;
	double TRNR8_p(t, z, y, x) ;
		TRNR8_p:long_name = "large particulate organic phosphorus" ;
		TRNR8_p:units = "mmol/m3" ;
	double TRNR8_s(t, z, y, x) ;
		TRNR8_s:long_name = "large particulate organic silicate" ;
		TRNR8_s:units = "mmol/m3" ;
	double TRNO2_o(t, z, y, x) ;
		TRNO2_o:long_name = "dissolved oxygen" ;
		TRNO2_o:units = "mmol/m3" ;
	double TRNO3_c(t, z, y, x) ;
		TRNO3_c:long_name = "dissolved inorganic carbon" ;
		TRNO3_c:units = "mmol/m3" ;
	double TRNO3_bioalk(t, z, y, x) ;
		TRNO3_bioalk:long_name = "biogeochemically induced alkalinity" ;
		TRNO3_bioalk:units = "umol/kg" ;
	double TRNN1_p(t, z, y, x) ;
		TRNN1_p:long_name = "phosphate" ;
		TRNN1_p:units = "mmol/m3" ;
	double TRNN3_n(t, z, y, x) ;
		TRNN3_n:long_name = "oxidised nitrogen" ;
		TRNN3_n:units = "mmol/m3" ;
	double TRNN4_n(t, z, y, x) ;
		TRNN4_n:long_name = "ammonium" ;
		TRNN4_n:units = "mmol/m3" ;
	double TRNN5_s(t, z, y, x) ;
		TRNN5_s:long_name = "silicate" ;
		TRNN5_s:units = "mmol/m3" ;
	double TRNL2_c(t, z, y, x) ;
		TRNL2_c:long_name = "calcite" ;
		TRNL2_c:units = "mg/m3" ;
	double TRNlight_ADY(t, z, y, x) ;
		TRNlight_ADY:long_name = "gelbstoff absoprtion" ;
		TRNlight_ADY:units = "1/m" ;
	double TRBP1_c(t, z, y, x) ;
		TRBP1_c:long_name = "diatom carbon" ;
		TRBP1_c:units = "mg/m3" ;
	double TRBP1_n(t, z, y, x) ;
		TRBP1_n:long_name = "diatom nitrogen" ;
		TRBP1_n:units = "mmol/m3" ;
	double TRBP1_p(t, z, y, x) ;
		TRBP1_p:long_name = "diatom phosphate" ;
		TRBP1_p:units = "mmol/m3" ;
	double TRBP1_s(t, z, y, x) ;
		TRBP1_s:long_name = "diatom silicate" ;
		TRBP1_s:units = "mmol/m3" ;
	double TRBP1_Chl(t, z, y, x) ;
		TRBP1_Chl:long_name = "diatom chlorophyll-a" ;
		TRBP1_Chl:units = "mg/m3" ;
	double TRBP2_c(t, z, y, x) ;
		TRBP2_c:long_name = "nanophytoplankton carbon" ;
		TRBP2_c:units = "mg/m3" ;
	double TRBP2_n(t, z, y, x) ;
		TRBP2_n:long_name = "nanophytoplankton nitrogen" ;
		TRBP2_n:units = "mmol/m3" ;
	double TRBP2_p(t, z, y, x) ;
		TRBP2_p:long_name = "nanophytoplankton phosphate" ;
		TRBP2_p:units = "mmol/m3" ;
	double TRBP2_Chl(t, z, y, x) ;
		TRBP2_Chl:long_name = "nanophytoplankton chlorophyll-a" ;
		TRBP2_Chl:units = "mg/m3" ;
	double TRBP3_c(t, z, y, x) ;
		TRBP3_c:long_name = "picophytoplankton carbon" ;
		TRBP3_c:units = "mg/m3" ;
	double TRBP3_n(t, z, y, x) ;
		TRBP3_n:long_name = "picophytoplankton nitrogen" ;
		TRBP3_n:units = "mmol/m3" ;
	double TRBP3_p(t, z, y, x) ;
		TRBP3_p:long_name = "picophytoplankton phosphate" ;
		TRBP3_p:units = "mmol/m3" ;
	double TRBP3_Chl(t, z, y, x) ;
		TRBP3_Chl:long_name = "picophytoplankton chlorophyll-a" ;
		TRBP3_Chl:units = "mg/m3" ;
	double TRBP4_c(t, z, y, x) ;
		TRBP4_c:long_name = "microphytoplankton carbon" ;
		TRBP4_c:units = "mg/m3" ;
	double TRBP4_n(t, z, y, x) ;
		TRBP4_n:long_name = "microphytoplankton nitrogen" ;
		TRBP4_n:units = "mmol/m3" ;
	double TRBP4_p(t, z, y, x) ;
		TRBP4_p:long_name = "microphytoplankton phosphate" ;
		TRBP4_p:units = "mmol/m3" ;
	double TRBP4_Chl(t, z, y, x) ;
		TRBP4_Chl:long_name = "microphytoplankton chlorophyll-a" ;
		TRBP4_Chl:units = "mg/m3" ;
	double TRBZ4_c(t, z, y, x) ;
		TRBZ4_c:long_name = "mesozooplankton carbon" ;
		TRBZ4_c:units = "mg/m3" ;
	double TRBZ5_c(t, z, y, x) ;
		TRBZ5_c:long_name = "microzooplankton carbon" ;
		TRBZ5_c:units = "mg/m3" ;
	double TRBZ5_n(t, z, y, x) ;
		TRBZ5_n:long_name = "microzooplankton nitrogen" ;
		TRBZ5_n:units = "mmol/m3" ;
	double TRBZ5_p(t, z, y, x) ;
		TRBZ5_p:long_name = "microzooplankton phosphorus" ;
		TRBZ5_p:units = "mmol/m3" ;
	double TRBZ6_c(t, z, y, x) ;
		TRBZ6_c:long_name = "heteroflagellates carbon" ;
		TRBZ6_c:units = "mg/m3" ;
	double TRBZ6_n(t, z, y, x) ;
		TRBZ6_n:long_name = "heteroflagellates nitrogen" ;
		TRBZ6_n:units = "mmol/m3" ;
	double TRBZ6_p(t, z, y, x) ;
		TRBZ6_p:long_name = "heteroflagellates phosphorus" ;
		TRBZ6_p:units = "mmol/m3" ;
	double TRBB1_c(t, z, y, x) ;
		TRBB1_c:long_name = "particualte organic carbon" ;
		TRBB1_c:units = "mg/m3" ;
	double TRBB1_n(t, z, y, x) ;
		TRBB1_n:long_name = "particualte organic nitrogen" ;
		TRBB1_n:units = "mmol/m3" ;
	double TRBB1_p(t, z, y, x) ;
		TRBB1_p:long_name = "particualte organic phosphorus" ;
		TRBB1_p:units = "mmol/m3" ;
	double TRBR1_c(t, z, y, x) ;
		TRBR1_c:long_name = "dissolved organic carbon" ;
		TRBR1_c:units = "mg/m3" ;
	double TRBR1_n(t, z, y, x) ;
		TRBR1_n:long_name = "dissolved organic nitrogen" ;
		TRBR1_n:units = "mmol/m3" ;
	double TRBR1_p(t, z, y, x) ;
		TRBR1_p:long_name = "dissolved organic phosphorus" ;
		TRBR1_p:units = "mmol/m3" ;
	double TRBR2_c(t, z, y, x) ;
		TRBR2_c:long_name = "semi-labile organic carbon" ;
		TRBR2_c:units = "mg/m3" ;
	double TRBR3_c(t, z, y, x) ;
		TRBR3_c:long_name = "semi-refractory organic carbon" ;
		TRBR3_c:units = "mg/m3" ;
	double TRBR4_c(t, z, y, x) ;
		TRBR4_c:long_name = "small particulate organic carbon" ;
		TRBR4_c:units = "mg/m3" ;
	double TRBR4_n(t, z, y, x) ;
		TRBR4_n:long_name = "small particulate organic nitrogen" ;
		TRBR4_n:units = "mmol/m3" ;
	double TRBR4_p(t, z, y, x) ;
		TRBR4_p:long_name = "small particulate organic phosphorus" ;
		TRBR4_p:units = "mmol/m3" ;
	double TRBR6_c(t, z, y, x) ;
		TRBR6_c:long_name = "medium size particulate organic carbon" ;
		TRBR6_c:units = "mg/m3" ;
	double TRBR6_n(t, z, y, x) ;
		TRBR6_n:long_name = "medium size particulate organic nitrogen" ;
		TRBR6_n:units = "mmol/m3" ;
	double TRBR6_p(t, z, y, x) ;
		TRBR6_p:long_name = "medium size particulate organic phosphorus" ;
		TRBR6_p:units = "mmol/m3" ;
	double TRBR6_s(t, z, y, x) ;
		TRBR6_s:long_name = "medium size particulate organic silicate" ;
		TRBR6_s:units = "mmol/m3" ;
	double TRBR8_c(t, z, y, x) ;
		TRBR8_c:long_name = "large particulate organic carbon" ;
		TRBR8_c:units = "mg/m3" ;
	double TRBR8_n(t, z, y, x) ;
		TRBR8_n:long_name = "large particulate organic nitrogen" ;
		TRBR8_n:units = "mmol/m3" ;
	double TRBR8_p(t, z, y, x) ;
		TRBR8_p:long_name = "large particulate organic phosphorus" ;
		TRBR8_p:units = "mmol/m3" ;
	double TRBR8_s(t, z, y, x) ;
		TRBR8_s:long_name = "large particulate organic silicate" ;
		TRBR8_s:units = "mmol/m3" ;
	double TRBO2_o(t, z, y, x) ;
		TRBO2_o:long_name = "dissolved oxygen" ;
		TRBO2_o:units = "mmol/m3" ;
	double TRBO3_c(t, z, y, x) ;
		TRBO3_c:long_name = "dissolved inorganic carbon" ;
		TRBO3_c:units = "mmol/m3" ;
	double TRBO3_bioalk(t, z, y, x) ;
		TRBO3_bioalk:long_name = "biogeochemically induced alkalinity" ;
		TRBO3_bioalk:units = "umol/kg" ;
	double TRBN1_p(t, z, y, x) ;
		TRBN1_p:long_name = "phosphate" ;
		TRBN1_p:units = "mmol/m3" ;
	double TRBN3_n(t, z, y, x) ;
		TRBN3_n:long_name = "oxidised nitrogen" ;
		TRBN3_n:units = "mmol/m3" ;
	double TRBN4_n(t, z, y, x) ;
		TRBN4_n:long_name = "ammonium" ;
		TRBN4_n:units = "mmol/m3" ;
	double TRBN5_s(t, z, y, x) ;
		TRBN5_s:long_name = "silicate" ;
		TRBN5_s:units = "mmol/m3" ;
	double TRBL2_c(t, z, y, x) ;
		TRBL2_c:long_name = "calcite" ;
		TRBL2_c:units = "mg/m3" ;
	double TRBlight_ADY(t, z, y, x) ;
		TRBlight_ADY:long_name = "gelbstoff absoprtion" ;
		TRBlight_ADY:units = "1/m" ;
	double fabm_st2DnH1_c(t, y, x) ;
		fabm_st2DnH1_c:long_name = "benthic aerobic bacteria" ;
		fabm_st2DnH1_c:units = "mmol/m2" ;
	double fabm_st2DnH2_c(t, y, x) ;
		fabm_st2DnH2_c:long_name = "benthic anaerobic bacteria" ;
		fabm_st2DnH2_c:units = "mmol/m2" ;
	double fabm_st2DnY2_c(t, y, x) ;
		fabm_st2DnY2_c:long_name = "deposit feeders" ;
		fabm_st2DnY2_c:units = "mg/m2" ;
	double fabm_st2DnY3_c(t, y, x) ;
		fabm_st2DnY3_c:long_name = "suspension feeders" ;
		fabm_st2DnY3_c:units = "mg/m2" ;
	double fabm_st2DnY4_c(t, y, x) ;
		fabm_st2DnY4_c:long_name = "meiobenthos" ;
		fabm_st2DnY4_c:units = "mg/m2" ;
	double fabm_st2DnQ1_c(t, y, x) ;
		fabm_st2DnQ1_c:long_name = "benthic dissolved organic carbon" ;
		fabm_st2DnQ1_c:units = "mg/m2" ;
	double fabm_st2DnQ1_n(t, y, x) ;
		fabm_st2DnQ1_n:long_name = "benthic dissolved organic nitrogen" ;
		fabm_st2DnQ1_n:units = "mmol/m2" ;
	double fabm_st2DnQ1_p(t, y, x) ;
		fabm_st2DnQ1_p:long_name = "benthic dissolved organic phosphorus" ;
		fabm_st2DnQ1_p:units = "mmol/m2" ;
	double fabm_st2DnQ6_c(t, y, x) ;
		fabm_st2DnQ6_c:long_name = "benthic particulate organic carbon" ;
		fabm_st2DnQ6_c:units = "mg/m2" ;
	double fabm_st2DnQ6_n(t, y, x) ;
		fabm_st2DnQ6_n:long_name = "benthic particulate organic nitrogen" ;
		fabm_st2DnQ6_n:units = "mmol/m2" ;
	double fabm_st2DnQ6_p(t, y, x) ;
		fabm_st2DnQ6_p:long_name = "benthic particulate organic phosphorus" ;
		fabm_st2DnQ6_p:units = "mmol/m2" ;
	double fabm_st2DnQ6_s(t, y, x) ;
		fabm_st2DnQ6_s:long_name = "benthic particulate organic silicate" ;
		fabm_st2DnQ6_s:units = "mmol/m2" ;
	double fabm_st2DnQ6_pen_depth_n(t, y, x) ;
		fabm_st2DnQ6_pen_depth_n:long_name = "penetration depth of benthic degradable nitrogen" ;
		fabm_st2DnQ6_pen_depth_n:units = "m" ;
	double fabm_st2DnQ6_pen_depth_c(t, y, x) ;
		fabm_st2DnQ6_pen_depth_c:long_name = "penetration depth of benthic degradable carbon" ;
		fabm_st2DnQ6_pen_depth_c:units = "m" ;
	double fabm_st2DnQ6_pen_depth_p(t, y, x) ;
		fabm_st2DnQ6_pen_depth_p:long_name = "penetration depth of benthic degradable phosphorus" ;
		fabm_st2DnQ6_pen_depth_p:units = "m" ;
	double fabm_st2DnQ6_pen_depth_s(t, y, x) ;
		fabm_st2DnQ6_pen_depth_s:long_name = "penetration depth of benthic degradable silicate" ;
		fabm_st2DnQ6_pen_depth_s:units = "m" ;
	double fabm_st2DnQ7_c(t, y, x) ;
		fabm_st2DnQ7_c:long_name = "benthic refractory organic carbon" ;
		fabm_st2DnQ7_c:units = "mg/m2" ;
	double fabm_st2DnQ7_n(t, y, x) ;
		fabm_st2DnQ7_n:long_name = "benthic refractory organic nitrogen" ;
		fabm_st2DnQ7_n:units = "mmol/m2" ;
	double fabm_st2DnQ7_p(t, y, x) ;
		fabm_st2DnQ7_p:long_name = "benthic refractory organic phosphorus" ;
		fabm_st2DnQ7_p:units = "mmol/m2" ;
	double fabm_st2DnQ7_pen_depth_c(t, y, x) ;
		fabm_st2DnQ7_pen_depth_c:long_name = "penetration depth of benthic refractory carbon" ;
		fabm_st2DnQ7_pen_depth_c:units = "m" ;
	double fabm_st2DnQ7_pen_depth_n(t, y, x) ;
		fabm_st2DnQ7_pen_depth_n:long_name = "penetration depth of benthic refractory nitrogen" ;
		fabm_st2DnQ7_pen_depth_n:units = "m" ;
	double fabm_st2DnQ7_pen_depth_p(t, y, x) ;
		fabm_st2DnQ7_pen_depth_p:long_name = "penetration depth of benthic refractory phosphorus" ;
		fabm_st2DnQ7_pen_depth_p:units = "m" ;
	double fabm_st2DnQ17_n(t, y, x) ;
		fabm_st2DnQ17_n:long_name = "benthic buried organic nitrogen" ;
		fabm_st2DnQ17_n:units = "mmol/m2" ;
	double fabm_st2DnQ17_c(t, y, x) ;
		fabm_st2DnQ17_c:long_name = "benthic buried organic carbon" ;
		fabm_st2DnQ17_c:units = "mg/m2" ;
	double fabm_st2DnQ17_p(t, y, x) ;
		fabm_st2DnQ17_p:long_name = "benthic buried organic phosphorus" ;
		fabm_st2DnQ17_p:units = "mmol/m2" ;
	double fabm_st2DnG2_o(t, y, x) ;
		fabm_st2DnG2_o:long_name = "benthic dissolved oxygen above oxygenated layer" ;
		fabm_st2DnG2_o:units = "mmol/m2" ;
	double fabm_st2DnG2_o_deep(t, y, x) ;
		fabm_st2DnG2_o_deep:long_name = "benthic dissolved oxygen below oxygenated layer" ;
		fabm_st2DnG2_o_deep:units = "mmol/m2" ;
	double fabm_st2DnG3_c(t, y, x) ;
		fabm_st2DnG3_c:long_name = "benthic dissolved inorganic carbon" ;
		fabm_st2DnG3_c:units = "mmol/m2" ;
	double fabm_st2DnK1_p(t, y, x) ;
		fabm_st2DnK1_p:long_name = "benthic phosphorus" ;
		fabm_st2DnK1_p:units = "mmol/m2" ;
	double fabm_st2DnK3_n(t, y, x) ;
		fabm_st2DnK3_n:long_name = "benthic nitrogen" ;
		fabm_st2DnK3_n:units = "mmol/m2" ;
	double fabm_st2DnK4_n(t, y, x) ;
		fabm_st2DnK4_n:long_name = "benthic ammonium" ;
		fabm_st2DnK4_n:units = "mmol/m2" ;
	double fabm_st2DnK5_s(t, y, x) ;
		fabm_st2DnK5_s:long_name = "benthic silicate" ;
		fabm_st2DnK5_s:units = "mmol/m2" ;
	double fabm_st2DnbL2_c(t, y, x) ;
		fabm_st2DnbL2_c:long_name = "calcite" ;
		fabm_st2DnbL2_c:units = "mg/m2" ;
	double fabm_st2Dnben_col_D2m(t, y, x) ;
		fabm_st2Dnben_col_D2m:long_name = "oxidised nitrogen horizon" ;
		fabm_st2Dnben_col_D2m:units = "m" ;
	double fabm_st2Dnben_col_D1m(t, y, x) ;
		fabm_st2Dnben_col_D1m:long_name = "dissolved oxygen horizon" ;
		fabm_st2Dnben_col_D1m:units = "m" ;
	double fabm_st2Dnben_nit_G4n(t, y, x) ;
		fabm_st2Dnben_nit_G4n:long_name = "benthic dinitrogen" ;
		fabm_st2Dnben_nit_G4n:units = "mmol/m2" ;
	double fabm_st2DbH1_c(t, y, x) ;
		fabm_st2DbH1_c:long_name = "benthic aerobic bacteria" ;
		fabm_st2DbH1_c:units = "mmol/m2" ;
	double fabm_st2DbH2_c(t, y, x) ;
		fabm_st2DbH2_c:long_name = "benthic anaerobic bacteria" ;
		fabm_st2DbH2_c:units = "mmol/m2" ;
	double fabm_st2DbY2_c(t, y, x) ;
		fabm_st2DbY2_c:long_name = "deposit feeders" ;
		fabm_st2DbY2_c:units = "mg/m2" ;
	double fabm_st2DbY3_c(t, y, x) ;
		fabm_st2DbY3_c:long_name = "suspension feeders" ;
		fabm_st2DbY3_c:units = "mg/m2" ;
	double fabm_st2DbY4_c(t, y, x) ;
		fabm_st2DbY4_c:long_name = "meiobenthos" ;
		fabm_st2DbY4_c:units = "mg/m2" ;
	double fabm_st2DbQ1_c(t, y, x) ;
		fabm_st2DbQ1_c:long_name = "benthic dissolved organic carbon" ;
		fabm_st2DbQ1_c:units = "mg/m2" ;
	double fabm_st2DbQ1_n(t, y, x) ;
		fabm_st2DbQ1_n:long_name = "benthic dissolved organic nitrogen" ;
		fabm_st2DbQ1_n:units = "mmol/m2" ;
	double fabm_st2DbQ1_p(t, y, x) ;
		fabm_st2DbQ1_p:long_name = "benthic dissolved organic phosphorus" ;
		fabm_st2DbQ1_p:units = "mmol/m2" ;
	double fabm_st2DbQ6_c(t, y, x) ;
		fabm_st2DbQ6_c:long_name = "benthic particulate organic carbon" ;
		fabm_st2DbQ6_c:units = "mg/m2" ;
	double fabm_st2DbQ6_n(t, y, x) ;
		fabm_st2DbQ6_n:long_name = "benthic particulate organic nitrogen" ;
		fabm_st2DbQ6_n:units = "mmol/m2" ;
	double fabm_st2DbQ6_p(t, y, x) ;
		fabm_st2DbQ6_p:long_name = "benthic particulate organic phosphorus" ;
		fabm_st2DbQ6_p:units = "mmol/m2" ;
	double fabm_st2DbQ6_s(t, y, x) ;
		fabm_st2DbQ6_s:long_name = "benthic particulate organic silicate" ;
		fabm_st2DbQ6_s:units = "mmol/m2" ;
	double fabm_st2DbQ6_pen_depth_n(t, y, x) ;
		fabm_st2DbQ6_pen_depth_n:long_name = "penetration depth of benthic degradable nitrogen" ;
		fabm_st2DbQ6_pen_depth_n:units = "m" ;
	double fabm_st2DbQ6_pen_depth_c(t, y, x) ;
		fabm_st2DbQ6_pen_depth_c:long_name = "penetration depth of benthic degradable carbon" ;
		fabm_st2DbQ6_pen_depth_c:units = "m" ;
	double fabm_st2DbQ6_pen_depth_p(t, y, x) ;
		fabm_st2DbQ6_pen_depth_p:long_name = "penetration depth of benthic degradable phosphorus" ;
		fabm_st2DbQ6_pen_depth_p:units = "m" ;
	double fabm_st2DbQ6_pen_depth_s(t, y, x) ;
		fabm_st2DbQ6_pen_depth_s:long_name = "penetration depth of benthic degradable silicate" ;
		fabm_st2DbQ6_pen_depth_s:units = "m" ;
	double fabm_st2DbQ7_c(t, y, x) ;
		fabm_st2DbQ7_c:long_name = "benthic refractory organic carbon" ;
		fabm_st2DbQ7_c:units = "mg/m2" ;
	double fabm_st2DbQ7_n(t, y, x) ;
		fabm_st2DbQ7_n:long_name = "benthic refractory organic nitrogen" ;
		fabm_st2DbQ7_n:units = "mmol/m2" ;
	double fabm_st2DbQ7_p(t, y, x) ;
		fabm_st2DbQ7_p:long_name = "benthic refractory organic phosphorus" ;
		fabm_st2DbQ7_p:units = "mmol/m2" ;
	double fabm_st2DbQ7_pen_depth_c(t, y, x) ;
		fabm_st2DbQ7_pen_depth_c:long_name = "penetration depth of benthic refractory carbon" ;
		fabm_st2DbQ7_pen_depth_c:units = "m" ;
	double fabm_st2DbQ7_pen_depth_n(t, y, x) ;
		fabm_st2DbQ7_pen_depth_n:long_name = "penetration depth of benthic refractory nitrogen" ;
		fabm_st2DbQ7_pen_depth_n:units = "m" ;
	double fabm_st2DbQ7_pen_depth_p(t, y, x) ;
		fabm_st2DbQ7_pen_depth_p:long_name = "penetration depth of benthic refractory phosphorus" ;
		fabm_st2DbQ7_pen_depth_p:units = "m" ;
	double fabm_st2DbQ17_n(t, y, x) ;
		fabm_st2DbQ17_n:long_name = "benthic buried organic nitrogen" ;
		fabm_st2DbQ17_n:units = "mmol/m2" ;
	double fabm_st2DbQ17_c(t, y, x) ;
		fabm_st2DbQ17_c:long_name = "benthic buried organic carbon" ;
		fabm_st2DbQ17_c:units = "mg/m2" ;
	double fabm_st2DbQ17_p(t, y, x) ;
		fabm_st2DbQ17_p:long_name = "benthic buried organic phosphorus" ;
		fabm_st2DbQ17_p:units = "mmol/m2" ;
	double fabm_st2DbG2_o(t, y, x) ;
		fabm_st2DbG2_o:long_name = "benthic dissolved oxygen above oxygenated layer" ;
		fabm_st2DbG2_o:units = "mmol/m2" ;
	double fabm_st2DbG2_o_deep(t, y, x) ;
		fabm_st2DbG2_o_deep:long_name = "benthic dissolved oxygen below oxygenated layer" ;
		fabm_st2DbG2_o_deep:units = "mmol/m2" ;
	double fabm_st2DbG3_c(t, y, x) ;
		fabm_st2DbG3_c:long_name = "benthic dissolved inorganic carbon" ;
		fabm_st2DbG3_c:units = "mmol/m2" ;
	double fabm_st2DbK1_p(t, y, x) ;
		fabm_st2DbK1_p:long_name = "benthic phosphorus" ;
		fabm_st2DbK1_p:units = "mmol/m2" ;
	double fabm_st2DbK3_n(t, y, x) ;
		fabm_st2DbK3_n:long_name = "benthic nitrogen" ;
		fabm_st2DbK3_n:units = "mmol/m2" ;
	double fabm_st2DbK4_n(t, y, x) ;
		fabm_st2DbK4_n:long_name = "benthic ammonium" ;
		fabm_st2DbK4_n:units = "mmol/m2" ;
	double fabm_st2DbK5_s(t, y, x) ;
		fabm_st2DbK5_s:long_name = "benthic silicate" ;
		fabm_st2DbK5_s:units = "mmol/m2" ;
	double fabm_st2DbbL2_c(t, y, x) ;
		fabm_st2DbbL2_c:long_name = "calcite" ;
		fabm_st2DbbL2_c:units = "mg/m2" ;
	double fabm_st2Dbben_col_D2m(t, y, x) ;
		fabm_st2Dbben_col_D2m:long_name = "oxidised nitrogen horizon" ;
		fabm_st2Dbben_col_D2m:units = "m" ;
	double fabm_st2Dbben_col_D1m(t, y, x) ;
		fabm_st2Dbben_col_D1m:long_name = "dissolved oxygen horizon" ;
		fabm_st2Dbben_col_D1m:units = "m" ;
	double fabm_st2Dbben_nit_G4n(t, y, x) ;
		fabm_st2Dbben_nit_G4n:long_name = "benthic dinitrogen" ;
		fabm_st2Dbben_nit_G4n:units = "mmol/m2" ;
}
